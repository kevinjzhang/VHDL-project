----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 13.10.2018 17:07:37
-- Design Name: 
-- Module Name: manchester_encoder_unit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity manchester_encoder_unit is
Port (hamming: in std_logic;
    manchester:out std_logic_vector(1 downto 0)
    );
end manchester_encoder_unit;

architecture Behavioral of manchester_encoder_unit is
    
begin
    manchester_dec: process(hamming)
    begin
        if hamming = '0' then
            manchester <= "10";
        else
            manchester <= "01";
        end if;
    end process;
end Behavioral;
